// copy queue contents to dynamic array
//1) I want to copy queue 1 into dynamic array and print it
//2) I want to copy dynmaic array into another queue 2
//3) Then copy queue 2 partially to queue 3 and print it
