// 1. Implement class based stack in SV
// 2. Extend the stack base class to implement FIFO
// 3. test your code and verify stack and fifo behaviour
